module top_module( 
    input [2:0] a,
    input [2:0] b,
    output [2:0] out_or_bitwise,
    output out_or_logical,
    output [5:0] out_not
);
    assign out_or_bitwise = a | b; // performs indipendent or operations of all bits 
    assign out_or_logical = a||b; // acts as a boolean function
    assign out_not[5:3] = ~b[2:0]; // inverses the bits of b
    assign out_not[2:0] = ~a[2:0]; // inverses the bits of a
endmodule
